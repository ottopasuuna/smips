`define AND    4'b0000
`define OR     4'b0001
`define ADD    4'b0010
`define SUB    4'b0110
`define SET_LT 4'b0111
`define NOR    4'b1100

