`define R_FORMAT 6'b000000
`define LW 6'b100011
`define SW 6'b101011
`define BEQ 6'b000100

